// de0_nano_system.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module de0_nano_system (
		output wire        clk100m_clk_clk,                           //                  clk100m_clk.clk
		input  wire        clk_50,                                    //                clk_50_clk_in.clk
		input  wire        reset_n,                                   //          clk_50_clk_in_reset.reset_n
		input  wire [1:0]  in_port_to_the_key,                        //      key_external_connection.export
		output wire [12:0] zs_addr_from_the_sdram,                    //                   sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                      //                             .ba
		output wire        zs_cas_n_from_the_sdram,                   //                             .cas_n
		output wire        zs_cke_from_the_sdram,                     //                             .cke
		output wire        zs_cs_n_from_the_sdram,                    //                             .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram,               //                             .dq
		output wire [1:0]  zs_dqm_from_the_sdram,                     //                             .dqm
		output wire        zs_ras_n_from_the_sdram,                   //                             .ras_n
		output wire        zs_we_n_from_the_sdram,                    //                             .we_n
		input  wire [3:0]  in_port_to_the_sw,                         //       sw_external_connection.export
		input  wire        trg_pls_component_0_spi_clk_clk,           //  trg_pls_component_0_spi_clk.clk
		input  wire        trg_pls_component_0_spi_cs_spi,            //   trg_pls_component_0_spi_cs.spi
		input  wire        trg_pls_component_0_spi_mosi_spi,          // trg_pls_component_0_spi_mosi.spi
		output wire [4:0]  trg_pls_component_0_trg_pls_triggersignal  //  trg_pls_component_0_trg_pls.triggersignal
	);

	wire         altpll_0_c1_clk;                                           // altpll_0:c1 -> TRG_PLS_component_0:CLK160M
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;             // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;              // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                 // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;            // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_trg_pls_component_0_reg_chipselect;      // mm_interconnect_0:TRG_PLS_component_0_reg_chipselect -> TRG_PLS_component_0:REG_CS
	wire  [31:0] mm_interconnect_0_trg_pls_component_0_reg_readdata;        // TRG_PLS_component_0:REG_READDATA -> mm_interconnect_0:TRG_PLS_component_0_reg_readdata
	wire         mm_interconnect_0_trg_pls_component_0_reg_waitrequest;     // TRG_PLS_component_0:REG_WAITREQUEST -> mm_interconnect_0:TRG_PLS_component_0_reg_waitrequest
	wire  [15:0] mm_interconnect_0_trg_pls_component_0_reg_address;         // mm_interconnect_0:TRG_PLS_component_0_reg_address -> TRG_PLS_component_0:REG_ADDRESS
	wire         mm_interconnect_0_trg_pls_component_0_reg_read;            // mm_interconnect_0:TRG_PLS_component_0_reg_read -> TRG_PLS_component_0:REG_READ
	wire         mm_interconnect_0_trg_pls_component_0_reg_begintransfer;   // mm_interconnect_0:TRG_PLS_component_0_reg_begintransfer -> TRG_PLS_component_0:REG_BEGINTRANSFER
	wire         mm_interconnect_0_trg_pls_component_0_reg_write;           // mm_interconnect_0:TRG_PLS_component_0_reg_write -> TRG_PLS_component_0:REG_WRITE
	wire  [31:0] mm_interconnect_0_trg_pls_component_0_reg_writedata;       // mm_interconnect_0:TRG_PLS_component_0_reg_writedata -> TRG_PLS_component_0:REG_WRITEDATA
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_key_s1_chipselect;                       // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                         // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                          // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_key_s1_write;                            // mm_interconnect_0:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                        // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire         mm_interconnect_0_sw_s1_chipselect;                        // mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                           // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_sw_s1_write;                             // mm_interconnect_0:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                         // mm_interconnect_0:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // key:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // sw:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller_001:reset_in0, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [jtag_uart:rst_n, key:reset_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, sdram:reset_n, sw:reset_n, timer:reset_n]
	wire         rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> [mm_interconnect_0:TRG_PLS_component_0_reg_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:TRG_PLS_component_0_reset_reset_bridge_in_reset_reset]

	ptmch_top trg_pls_component_0 (
		.RESET_N           (reset_n),                                                 //    reset.reset_n
		.REG_BEGINTRANSFER (mm_interconnect_0_trg_pls_component_0_reg_begintransfer), //      reg.begintransfer
		.REG_ADDRESS       (mm_interconnect_0_trg_pls_component_0_reg_address),       //         .address
		.REG_READ          (mm_interconnect_0_trg_pls_component_0_reg_read),          //         .read
		.REG_WRITE         (mm_interconnect_0_trg_pls_component_0_reg_write),         //         .write
		.REG_READDATA      (mm_interconnect_0_trg_pls_component_0_reg_readdata),      //         .readdata
		.REG_WRITEDATA     (mm_interconnect_0_trg_pls_component_0_reg_writedata),     //         .writedata
		.REG_WAITREQUEST   (mm_interconnect_0_trg_pls_component_0_reg_waitrequest),   //         .waitrequest
		.REG_CS            (mm_interconnect_0_trg_pls_component_0_reg_chipselect),    //         .chipselect
		.CLK100M           (clk100m_clk_clk),                                         //  CLK100M.clk
		.CLK160M           (altpll_0_c1_clk),                                         //  CLK160M.clk
		.SPI_CLK           (trg_pls_component_0_spi_clk_clk),                         //  SPI_CLK.clk
		.SPI_CS            (trg_pls_component_0_spi_cs_spi),                          //   SPI_CS.spi
		.SPI_MOSI          (trg_pls_component_0_spi_mosi_spi),                        // SPI_MOSI.spi
		.TRG_PLS           (trg_pls_component_0_trg_pls_triggersignal)                //  TRG_PLS.triggersignal
	);

	de0_nano_system_altpll_0 altpll_0 (
		.clk                (clk_50),                                         //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (clk100m_clk_clk),                                //                    c0.clk
		.c1                 (altpll_0_c1_clk),                                //                    c1.clk
		.areset             (),                                               //        areset_conduit.export
		.locked             (),                                               //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	de0_nano_system_cpu cpu (
		.clk                                 (clk100m_clk_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	de0_nano_system_jtag_uart jtag_uart (
		.clk            (clk100m_clk_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	de0_nano_system_key key (
		.clk        (clk100m_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_key),                  // external_connection.export
		.irq        (irq_mapper_receiver1_irq)             //                 irq.irq
	);

	de0_nano_system_sdram sdram (
		.clk            (clk100m_clk_clk),                          //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	de0_nano_system_sw sw (
		.clk        (clk100m_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),    //                    .readdata
		.in_port    (in_port_to_the_sw),                   // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	de0_nano_system_timer timer (
		.clk        (clk100m_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	de0_nano_system_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                                      (clk100m_clk_clk),                                           //                                                    altpll_0_c0.clk
		.clk_50_clk_clk                                                       (clk_50),                                                    //                                                     clk_50_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                            //           altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                                (rst_controller_001_reset_out_reset),                        //                                cpu_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset                          (rst_controller_002_reset_out_reset),                        //                          jtag_uart_reset_reset_bridge_in_reset.reset
		.TRG_PLS_component_0_reg_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                        // TRG_PLS_component_0_reg_translator_reset_reset_bridge_in_reset.reset
		.TRG_PLS_component_0_reset_reset_bridge_in_reset_reset                (rst_controller_003_reset_out_reset),                        //                TRG_PLS_component_0_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                              (cpu_data_master_address),                                   //                                                cpu_data_master.address
		.cpu_data_master_waitrequest                                          (cpu_data_master_waitrequest),                               //                                                               .waitrequest
		.cpu_data_master_byteenable                                           (cpu_data_master_byteenable),                                //                                                               .byteenable
		.cpu_data_master_read                                                 (cpu_data_master_read),                                      //                                                               .read
		.cpu_data_master_readdata                                             (cpu_data_master_readdata),                                  //                                                               .readdata
		.cpu_data_master_write                                                (cpu_data_master_write),                                     //                                                               .write
		.cpu_data_master_writedata                                            (cpu_data_master_writedata),                                 //                                                               .writedata
		.cpu_data_master_debugaccess                                          (cpu_data_master_debugaccess),                               //                                                               .debugaccess
		.cpu_instruction_master_address                                       (cpu_instruction_master_address),                            //                                         cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                   (cpu_instruction_master_waitrequest),                        //                                                               .waitrequest
		.cpu_instruction_master_read                                          (cpu_instruction_master_read),                               //                                                               .read
		.cpu_instruction_master_readdata                                      (cpu_instruction_master_readdata),                           //                                                               .readdata
		.altpll_0_pll_slave_address                                           (mm_interconnect_0_altpll_0_pll_slave_address),              //                                             altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                             (mm_interconnect_0_altpll_0_pll_slave_write),                //                                                               .write
		.altpll_0_pll_slave_read                                              (mm_interconnect_0_altpll_0_pll_slave_read),                 //                                                               .read
		.altpll_0_pll_slave_readdata                                          (mm_interconnect_0_altpll_0_pll_slave_readdata),             //                                                               .readdata
		.altpll_0_pll_slave_writedata                                         (mm_interconnect_0_altpll_0_pll_slave_writedata),            //                                                               .writedata
		.cpu_debug_mem_slave_address                                          (mm_interconnect_0_cpu_debug_mem_slave_address),             //                                            cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                            (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                                               .write
		.cpu_debug_mem_slave_read                                             (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                                               .read
		.cpu_debug_mem_slave_readdata                                         (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                                               .readdata
		.cpu_debug_mem_slave_writedata                                        (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                                               .writedata
		.cpu_debug_mem_slave_byteenable                                       (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                                               .byteenable
		.cpu_debug_mem_slave_waitrequest                                      (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                                               .waitrequest
		.cpu_debug_mem_slave_debugaccess                                      (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                                               .debugaccess
		.jtag_uart_avalon_jtag_slave_address                                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                                    jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                               .write
		.jtag_uart_avalon_jtag_slave_read                                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                               .read
		.jtag_uart_avalon_jtag_slave_readdata                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                               .readdata
		.jtag_uart_avalon_jtag_slave_writedata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                               .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                               .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                               .chipselect
		.key_s1_address                                                       (mm_interconnect_0_key_s1_address),                          //                                                         key_s1.address
		.key_s1_write                                                         (mm_interconnect_0_key_s1_write),                            //                                                               .write
		.key_s1_readdata                                                      (mm_interconnect_0_key_s1_readdata),                         //                                                               .readdata
		.key_s1_writedata                                                     (mm_interconnect_0_key_s1_writedata),                        //                                                               .writedata
		.key_s1_chipselect                                                    (mm_interconnect_0_key_s1_chipselect),                       //                                                               .chipselect
		.sdram_s1_address                                                     (mm_interconnect_0_sdram_s1_address),                        //                                                       sdram_s1.address
		.sdram_s1_write                                                       (mm_interconnect_0_sdram_s1_write),                          //                                                               .write
		.sdram_s1_read                                                        (mm_interconnect_0_sdram_s1_read),                           //                                                               .read
		.sdram_s1_readdata                                                    (mm_interconnect_0_sdram_s1_readdata),                       //                                                               .readdata
		.sdram_s1_writedata                                                   (mm_interconnect_0_sdram_s1_writedata),                      //                                                               .writedata
		.sdram_s1_byteenable                                                  (mm_interconnect_0_sdram_s1_byteenable),                     //                                                               .byteenable
		.sdram_s1_readdatavalid                                               (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                                               .readdatavalid
		.sdram_s1_waitrequest                                                 (mm_interconnect_0_sdram_s1_waitrequest),                    //                                                               .waitrequest
		.sdram_s1_chipselect                                                  (mm_interconnect_0_sdram_s1_chipselect),                     //                                                               .chipselect
		.sw_s1_address                                                        (mm_interconnect_0_sw_s1_address),                           //                                                          sw_s1.address
		.sw_s1_write                                                          (mm_interconnect_0_sw_s1_write),                             //                                                               .write
		.sw_s1_readdata                                                       (mm_interconnect_0_sw_s1_readdata),                          //                                                               .readdata
		.sw_s1_writedata                                                      (mm_interconnect_0_sw_s1_writedata),                         //                                                               .writedata
		.sw_s1_chipselect                                                     (mm_interconnect_0_sw_s1_chipselect),                        //                                                               .chipselect
		.timer_s1_address                                                     (mm_interconnect_0_timer_s1_address),                        //                                                       timer_s1.address
		.timer_s1_write                                                       (mm_interconnect_0_timer_s1_write),                          //                                                               .write
		.timer_s1_readdata                                                    (mm_interconnect_0_timer_s1_readdata),                       //                                                               .readdata
		.timer_s1_writedata                                                   (mm_interconnect_0_timer_s1_writedata),                      //                                                               .writedata
		.timer_s1_chipselect                                                  (mm_interconnect_0_timer_s1_chipselect),                     //                                                               .chipselect
		.TRG_PLS_component_0_reg_address                                      (mm_interconnect_0_trg_pls_component_0_reg_address),         //                                        TRG_PLS_component_0_reg.address
		.TRG_PLS_component_0_reg_write                                        (mm_interconnect_0_trg_pls_component_0_reg_write),           //                                                               .write
		.TRG_PLS_component_0_reg_read                                         (mm_interconnect_0_trg_pls_component_0_reg_read),            //                                                               .read
		.TRG_PLS_component_0_reg_readdata                                     (mm_interconnect_0_trg_pls_component_0_reg_readdata),        //                                                               .readdata
		.TRG_PLS_component_0_reg_writedata                                    (mm_interconnect_0_trg_pls_component_0_reg_writedata),       //                                                               .writedata
		.TRG_PLS_component_0_reg_begintransfer                                (mm_interconnect_0_trg_pls_component_0_reg_begintransfer),   //                                                               .begintransfer
		.TRG_PLS_component_0_reg_waitrequest                                  (mm_interconnect_0_trg_pls_component_0_reg_waitrequest),     //                                                               .waitrequest
		.TRG_PLS_component_0_reg_chipselect                                   (mm_interconnect_0_trg_pls_component_0_reg_chipselect)       //                                                               .chipselect
	);

	de0_nano_system_irq_mapper irq_mapper (
		.clk           (clk100m_clk_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                       // reset_in0.reset
		.clk            (clk_50),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (cpu_debug_reset_request_reset),          // reset_in0.reset
		.clk            (clk100m_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk100m_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (clk100m_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
