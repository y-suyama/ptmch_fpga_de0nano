//==================================================================================================
//  Company name        : 
//  Date                : 
//  File Name           : ptmch_top_tb.sv
//  Project Name        : 
//  Coding              : suyama
//  Rev.                : 1.0
//
//==================================================================================================
// time scale
//==================================================================================================
    `timescale 1ns/1ps
//==================================================================================================
// Module
//==================================================================================================
module ptmch_top_tb();
    // Reset/Clock
    logic         RESET_N;
    logic         CLK160M;
    logic         CLK100M;
    // SPI Interface
    logic         SPI_CS;
    logic         SPI_CLK;
    logic         SPI_MOSI;
    logic [ 4: 0] TRG_PLS;
    // Avalone Slave I/F
    logic         REG_BEGINTRANSFER;
    logic [12: 0] REG_ADDRESS;
    logic         REG_CS;
    logic         REG_READ;
    logic         REG_WRITE;
    logic [31: 0] REG_READDATA;
    logic [31: 0] REG_WRITEDATA;
    logic         REG_WAITREQUEST;

//==================================================================================================
//  Structural coding
//==================================================================================================
ptmch_top _ptmch_top(
    .RESET_N(RESET_N),
    .CLK160M(CLK160M),
    .CLK100M(CLK100M),
    .SPI_CS(SPI_CS),
    .SPI_CLK(SPI_CLK),
    .SPI_MOSI(SPI_MOSI),
    .TRG_PLS(TRG_PLS),
    .REG_BEGINTRANSFER(REG_BEGINTRANSFER),
    .REG_ADDRESS(REG_ADDRESS),
    .REG_CS(REG_CS),
    .REG_READ(REG_READ),
    .REG_WRITE(REG_WRITE),
    .REG_READDATA(REG_READDATA),
    .REG_WRITEDATA(REG_WRITEDATA),
    .REG_WAITREQUEST(REG_WAITREQUEST)
);
//==================================================================================================
//  PARAMETER declarations
//==================================================================================================
    parameter cycle_160m         = 6.25;
    parameter half_cycle_160m    = 3.125;
    parameter half_cycle_100m    = 5;
    parameter cycle_spi          = 10;
    parameter half_cycle_spi     = 5;
    parameter start_delay        = 100;
    parameter cs_delay           = 200;
    parameter clk_delay          = 300;
//==================================================================================================
//  RESET/Clock
//==================================================================================================
    // PLL Clock 100MHz
    always #half_cycle_100m CLK100M = ~CLK100M;
    // PLL Clock 200MHz
    always #half_cycle_160m CLK160M = ~CLK160M;
//==================================================================================================
//  Initial
//==================================================================================================
    initial begin

        RESET_N  = 1'b1;
        CLK160M  = 1'b1;
        CLK100M  = 1'b1;
        SPI_CS   = 1'b1;
        SPI_CLK  = 1'b0;
        SPI_MOSI = 1'b1;
        REG_BEGINTRANSFER = 1'b0;
        REG_ADDRESS = 13'b0;
        REG_CS = 1'b0;
        REG_READ = 1'b0;
        REG_WRITE = 1'b0;
        REG_READDATA = 32'b0;
        REG_WRITEDATA = 32'b0;
        REG_WAITREQUEST = 1'b0;

        #start_delay    RESET_N = 1'b0;
        #start_delay    RESET_N = 1'b1;
        // program_excute 1 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // program_excute 2 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b1;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // program_excute 3 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b1;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // readstatus 1 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // readstatus 2 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b1;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // readstatus 3 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // 128kb_blockerase 1 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b1;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // 128kb_blockerase 2 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // 128kb_blockerase 3 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b1;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // pagedata_read 1 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // pagedata_read 2 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // pagedata_read 3 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // writestatus1 1 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                         SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                       SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // pagedata_read 2 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
        // pagedata_read 3 time
        #cs_delay       SPI_CS = 1'b0;
        #clk_delay      SPI_MOSI = 1'b0;//[7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        // Page Address
                        SPI_MOSI = 1'b0;//[23]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[22]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[21]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[20]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[19]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[18]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[17]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[16]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[15]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[14]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[13]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[12]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[11]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[10]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 9]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 8]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 7]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 6]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 5]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 4]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 3]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 2]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b0;//[ 1]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_MOSI = 1'b1;//[ 0]
        #half_cycle_spi SPI_CLK = 1'b1;
        #half_cycle_spi SPI_CLK = 1'b0;
        #half_cycle_spi SPI_CLK = 1'b0;
                        SPI_CS = 1'b1;
//        $finish;
   end
endmodule
